package pkg_arbiter_types;

parameter CLK_PERIOD = 10;
parameter NUMUNITS = 8;
parameter ADDRESSWIDTH = 3; //number of bits needed to address NUMUNITS
parameter NB_TRANSACTION_GENERATED = 64;

endpackage : pkg_arbiter_types